`ifndef BUF_INSTRUCTIONS
    `define BUF_INSTRUCTIONS 1

    `define BUF_IDLE_TWO      0;
    `define BUF_LOAD_TWO      1; // Take from a BUS and keep
    `define BUF_STORE_TWO     2; // Put the register value on a BUS
`endif
