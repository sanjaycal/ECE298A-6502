`ifndef ALU_OPCODES

    `define ALU_OPCODES 1
    //OPCODE
    `define NOP 3'b000
    `define ASL 3'b001


`endif
