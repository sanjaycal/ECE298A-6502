`ifndef ALU_OPCODES

    `define ALU_OPCODES 1
    //OPCODE
    `define NOP 4'b0000
    `define ASL 4'b0001

    `define ADR 4'b1110
    `define TMX 4'b1111


`endif
