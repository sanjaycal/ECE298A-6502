`ifndef ALU_OPCODES

    `define ALU_OPCODES 1
    //OPCODE
    `define NOP 4'b0000
    `define ASL 4'b0001
    `define LSR 4'b0010

    `define ADD 4'b1110
    `define TMX 4'b1111


`endif
