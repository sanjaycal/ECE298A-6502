`ifndef ALU_OPCODES

    `define ALU_OPCODES 1
    //OPCODE
    `define NOP 5'b00000
    `define ASL 5'b00001
    `define LSR 5'b00010
    `define ROL 5'b00011
    `define ROR 5'b00100
    `define AND 5'b00101
    `define OR 5'b00110


    `define FLG 5'b11101
    `define ADD 5'b11110
    `define TMX 5'b11111


`endif
