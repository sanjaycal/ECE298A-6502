`ifndef OPCODES
    //OPCODE
    `define NOP 8'000
    `define ASL 8'001


`endif
